`include "errors_base_vseq.sv"

`include "power_loss_seq.sv"
`include "power_loss_vseq.sv"