`include "../user_sequences/user_base_seq.sv"

`include "../user_sequences/simple_test_seq.sv"
`include "../user_sequences/one_coin_seq.sv"
`include "../user_sequences/few_coin_seq.sv"
`include "../user_sequences/dollars_seq.sv"
`include "../user_sequences/euros_seq.sv"
`include "../user_sequences/random_client_with_no_change_seq.sv"
`include "../user_sequences/full_client_session_with_no_errors_seq.sv"
`include "../user_sequences/lots_of_purchases_seq.sv"

`include "../user_sequences/buy_one_item_seq.sv"