`ifndef USER_SEQUENCES_INC
`define USER_SEQUENCES_INC

    `include "../user_sequences/user_base_seq.sv"

    `include "../user_sequences/simple_test_seq.sv"
    `include "../user_sequences/test_one_coin_seq.sv"
    `include "../user_sequences/test_few_coin_seq.sv"
    `include "../user_sequences/test_dollars_seq.sv"
    `include "../user_sequences/test_euros_seq.sv"
    `include "../user_sequences/test_random_client_with_no_change_seq.sv"
    `include "../user_sequences/full_client_session_with_no_errors_seq.sv"
    `include "../user_sequences/test_lots_of_purchases_seq.sv"

    `include "../user_sequences/buy_one_product_seq.sv"

`endif