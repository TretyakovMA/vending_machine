`ifndef REGISTER_SEQUENCES_INC
`define REGISTER_SEQUENCES_INC

`include "base_reg_seq.sv"

`include "register_test_vseq.sv"
`include "read_after_reset_test_seq.sv"
`include "read_after_write_test_seq.sv"

`include "change_item_price_seq.sv"


`endif