`ifndef READ_AFTER_WRITE_TEST
`define READ_AFTER_WRITE_TEST
class read_after_write_test extends register_base_test #(
	read_after_write_test_seq
);
	`uvm_component_utils(read_after_write_test)
	
	function new(string name = "read_after_write_test", uvm_component parent);
		super.new(name, parent);
	endfunction
	
	
endclass
`endif