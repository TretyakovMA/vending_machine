`include "interfaces/user_interface.sv"
`include "interfaces/register_interface.sv"
`include "interfaces/errors_interface.sv"
`include "interfaces/admin_interface.sv"