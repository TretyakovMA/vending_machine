`include "../integration_sequences/integration_base_virtual_seq.sv"

`include "../integration_sequences/buy_one_item_after_change_price_vseq.sv"
`include "../integration_sequences/c_s_after_change_price_vseq.sv"
`include "../integration_sequences/c_s_after_change_discount_vseq.sv"
`include "../integration_sequences/c_s_after_change_exchange_rate_vseq.sv"
`include "../integration_sequences/c_s_after_change_all_registers_vseq.sv"  
`include "../integration_sequences/c_s_with_interrupt_vseq.sv"  