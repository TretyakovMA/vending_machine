`include "user_tests/user_base_test.sv"
//`include "user_tests/simple_test.sv"
//`include "user_tests/test_one_coin.sv"
//`include "user_tests/test_few_coin.sv"
//`include "user_tests/test_dollars.sv"
//`include "user_tests/test_euros.sv"
//`include "user_tests/test_random_client_with_no_change.sv"
//`include "user_tests/full_client_session_with_no_errors.sv"
`include "user_tests/test_lots_of_purchases.sv"