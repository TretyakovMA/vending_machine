`include "register_tests/register_base_test.sv"
`include "register_tests/register_test.sv"