`include "../emergency_sequences/activate_emergency_signals_seq.sv"