`include "user_interface.sv"
`include "register_interface.sv"
`include "errors_interface.sv"
`include "admin_interface.sv"