`include "register_sequences/base_reg_seq.sv"

`include "register_sequences/register_test_seq.sv"
`include "register_sequences/register_test_vseq.sv"