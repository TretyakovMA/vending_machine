`ifndef ENVIROMENT_INC
`define ENVIROMENT_INC

    `include "env_config.sv"
	`include "env.sv"
	`include "base_test.sv"
	`include "sequence_base_test.sv"

`endif