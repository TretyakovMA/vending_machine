`ifndef REGISTERS_INC
`define REGISTERS_INC

    `include "../registers/vend_cfg_reg.sv"
    `include "../registers/vend_clients_reg.sv"
    `include "../registers/vend_item_reg.sv"
    `include "../registers/vend_paswd_reg.sv"
    `include "../registers/vm_reg_block.sv"

`endif