`include "../error_sequences/activate_error_signals_seq.sv"