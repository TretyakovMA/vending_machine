`include "../admin_sequences/admin_mode_on_seq.sv"
`include "../admin_sequences/admin_mode_off_seq.sv"