`include "vm_scoreboard.sv"
`include "vm_coverage.sv"