`include "base_macros.svh"
`include "my_report_server.sv"

`include "void_monitor.sv"
`include "void_driver.sv"

`include "base_transaction.sv"
`include "base_agent_config.sv"
`include "base_driver.sv"
`include "base_monitor.sv"
	
`include "base_agent.sv"
