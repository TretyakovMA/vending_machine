`ifndef SUMMARY_TESTS_INC
`define SUMMARY_TESTS_INC

`include "summary_base_test.sv"

`include "buy_one_product_test.sv"
`include "client_session_after_write_reg_test.sv"

`endif