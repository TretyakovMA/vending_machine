`include "../error_tests/check_alarm_test.sv"