`include "register_base_test.sv"

`include "read_after_reset_test.sv"
`include "read_after_write_test.sv"