`include "../integration_tests/integration_base_test.sv"

`include "../integration_tests/buy_one_item_after_change_price_test.sv"
`include "../integration_tests/c_s_after_change_price_test.sv"
`include "../integration_tests/c_s_after_change_discount_test.sv"
`include "../integration_tests/c_s_after_change_exchange_rate_test.sv"
`include "../integration_tests/c_s_after_change_all_registers_test.sv"

`include "../integration_tests/c_s_with_emergency_test.sv"
`include "../integration_tests/write_registers_with_emergency_test.sv"

`include "../integration_tests/c_s_with_reset_test.sv"