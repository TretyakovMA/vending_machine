`include "errors_transaction.sv"
`include "errors_driver.sv"
typedef uvm_sequencer #(errors_transaction) errors_sequencer;
`include "errors_agent.sv"