`include "../register_sequences/register_base_seq.sv"
`include "../register_sequences/register_base_virtual_seq.sv"
    
`include "../register_sequences/check_after_reset_seq.sv"
`include "../register_sequences/check_write_seq.sv"
`include "../register_sequences/check_read_seq.sv"

`include "../register_sequences/change_item_price_seq.sv"
`include "../register_sequences/change_item_discount_seq.sv"
`include "../register_sequences/change_exchange_rate_seq.sv"
`include "../register_sequences/change_all_registers_seq.sv"

`include "../register_sequences/write_registers_with_emergency_seq.sv"