`include "user_interface.sv"
`include "admin_interface.sv"
`include "register_interface.sv"
`include "emergency_interface.sv"