`ifndef REGISTER_TESTS_INC
`define REGISTER_TESTS_INC

    `include "../register_tests/register_base_test.sv"

    `include "../register_tests/read_after_reset_test.sv"
    `include "../register_tests/read_after_write_test.sv"
    
`endif