`include "../emergency_tests/check_alarm_test.sv"