`include "../register_tests/register_base_test.sv"

`include "../register_tests/check_after_reset_test.sv"
`include "../register_tests/check_write_test.sv"
`include "../register_tests/check_read_test.sv"
