`include "errors_base_test.sv"

`include "power_loss_test.sv"