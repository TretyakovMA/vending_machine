`ifndef RESET_INTERFACE
`define RESET_INTERFACE
interface reset_interface (input clk);

    logic rst_n;
    
endinterface
`endif