`include "../reset_sequences/initial_reset_seq.sv"
`include "../reset_sequences/reset_seq.sv"