`include "../reset_sequences/initial_reset_seq.sv"
`include "../reset_sequences/activate_reset_seq.sv"