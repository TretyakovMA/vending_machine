`ifndef SUMMARY_TESTS_INC
`define SUMMARY_TESTS_INC

`include "summary_base_test.sv"

`include "buy_one_product_test.sv"

`endif