`ifndef SUMMARY_SEQUENCES_INC
`define SUMMARY_SEQUENCES_INC

`include "summary_base_vseq.sv"

`include "buy_one_product_vseq.sv"

`endif