`include "vm_base_driver.sv"
`include "vm_base_monitor.sv"