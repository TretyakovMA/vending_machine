`ifndef FULL_INTERFACE 
`define FULL_INTERFACE

    `include "user_interface.sv"
    `include "register_interface.sv"
    `include "errors_interface.sv"
    `include "admin_interface.sv"
    
`endif