`include "sequence_base_test.sv"
`include "env_config.sv"
`include "env.sv"
`include "initiator.sv"
`include "base_test.sv"