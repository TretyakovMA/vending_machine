`define NUM_ITEMS 10
`define MAX_CLIENTS 100

`include "interfaces/user_interface.sv"
`include "interfaces/register_interface.sv"
`include "interfaces/errors_interface.sv"
`include "interfaces/admin_interface.sv"